`timescale 1ns / 1ps


module aes
    #(
        parameter int unsigned STATE_ARRAY_SIZE
    )
    (
        input logic state_array[STATE_ARRAY_SIZE/2][STATE_ARRAY_SIZE/2]


    );



endmodule
